module GX4000_video
(
    input         clk_sys,
    input         reset,
    input         gx4000_mode,
    input         plus_mode,
    
    // CPU interface
    input  [15:0] cpu_addr,
    input   [7:0] cpu_data,
    input         cpu_wr,
    input         cpu_rd,
    
    // Video input
    input   [1:0] r_in,
    input   [1:0] g_in,
    input   [1:0] b_in,
    input         hblank,
    input         vblank,
    
    // Sprite interface
    input   [7:0] sprite_pixel,
    input         sprite_active,
    input   [3:0] sprite_id,
    
    // Video output
    output  [1:0] r_out,
    output  [1:0] g_out,
    output  [1:0] b_out,
    
    // Collision detection
    output  [7:0] collision_reg,
    
    // Configuration interface
    output  [7:0] config_reg
);

    // Color palette registers
    reg [23:0] palette[0:31]; // 32 colors, 24-bit RGB
    
    // Video registers
    reg [7:0] screen_x;
    reg [7:0] screen_y;
    reg [7:0] video_mode;
    reg [7:0] collision_flags;
    
    // Sprite transformation registers
    reg [7:0] sprite_scale_x[0:7];
    reg [7:0] sprite_scale_y[0:7];
    reg [7:0] sprite_rotation[0:7];
    reg [7:0] sprite_center_x[0:7];
    reg [7:0] sprite_center_y[0:7];
    reg [7:0] sprite_alpha[0:7];
    reg [7:0] sprite_flip_x[0:7];
    reg [7:0] sprite_flip_y[0:7];
    reg [7:0] sprite_priority[0:7];
    reg [7:0] sprite_effect[0:7];
    
    // Video state
    reg [1:0] r_reg;
    reg [1:0] g_reg;
    reg [1:0] b_reg;
    reg [2:0] active_sprite;
    
    // Configuration registers
    reg [7:0] config_mode;
    reg [7:0] config_palette;
    reg [7:0] config_sprite;
    reg [7:0] config_video;
    reg [7:0] config_audio;
    reg [7:0] config_io;
    
    // Configuration presets
    reg [7:0] config_preset;
    reg [7:0] config_save[0:7];
    reg [7:0] config_load[0:7];
    
    // Previous color registers for effects
    reg [7:0] r_reg_prev;
    reg [7:0] g_reg_prev;
    reg [7:0] b_reg_prev;
    
    // Frame counter for effects
    reg [7:0] frame_counter;
    
    // Sprite transformation registers
    reg [7:0] angle;
    reg [7:0] scale_x;
    reg [7:0] scale_y;
    reg [7:0] center_x;
    reg [7:0] center_y;
    
    // Rotation registers
    reg [15:0] cos_angle;
    reg [15:0] sin_angle;
    reg [15:0] rot_x;
    reg [15:0] rot_y;
    
    // Position registers
    reg [7:0] final_x;
    reg [7:0] final_y;
    
    // Video effect registers
    reg [7:0] gray;
    reg [7:0] wave_offset;
    reg [7:0] wave_x;
    reg [7:0] zoom_x;
    reg [7:0] zoom_y;
    reg [7:0] cycle_offset;
    
    // Alpha blending registers
    logic [7:0] alpha;
    
    // Sine/Cosine lookup table for sprite rotation
    reg [7:0] sin_table[0:255];
    reg [7:0] cos_table[0:255];
    
    // Initialize lookup tables with pre-calculated fixed-point values
    initial begin
        // Pre-calculated sine values (scaled to 8-bit signed)
        for (int i = 0; i < 256; i = i + 1) begin
            // Convert angle to radians and calculate sin/cos
            // Scale to 8-bit signed value (-128 to 127)
            // Use fixed-point arithmetic instead of $rtoi
            sin_table[i] = (i < 128) ? (i * 127 / 128) : ((256 - i) * 127 / 128);
            cos_table[i] = (i < 64) ? (127 - (i * 127 / 64)) : 
                          (i < 192) ? ((i - 64) * 127 / 128 - 127) : 
                          (127 - ((i - 192) * 127 / 64));
        end
    end
    
    // Video processing
    always @(posedge clk_sys) begin
        if (reset) begin
            for (integer i = 0; i < 32; i = i + 1) begin
                palette[i] <= 24'h000000;
            end
            screen_x <= 8'h00;
            screen_y <= 8'h00;
            video_mode <= 8'h00;
            collision_flags <= 8'h00;
            r_reg <= 2'h0;
            g_reg <= 2'h0;
            b_reg <= 2'h0;
            active_sprite <= 3'h0;
            
            // Initialize sprite transformations
            for (integer i = 0; i < 8; i = i + 1) begin
                sprite_scale_x[i] <= 8'h40; // 1.0 scale
                sprite_scale_y[i] <= 8'h40; // 1.0 scale
                sprite_rotation[i] <= 8'h00; // 0 degrees
                sprite_center_x[i] <= 8'h00;
                sprite_center_y[i] <= 8'h00;
                sprite_alpha[i] <= 8'hFF; // Fully opaque
                sprite_flip_x[i] <= 8'h00;
                sprite_flip_y[i] <= 8'h00;
                sprite_priority[i] <= 8'h00;
                sprite_effect[i] <= 8'h00;
            end
            
            // Initialize configuration
            config_mode <= 8'h00;
            config_palette <= 8'h00;
            config_sprite <= 8'h00;
            config_video <= 8'h00;
            config_audio <= 8'h00;
            config_io <= 8'h00;
            config_preset <= 8'h00;
            
            // Initialize presets
            for (integer i = 0; i < 8; i = i + 1) begin
                config_save[i] <= 8'h00;
                config_load[i] <= 8'h00;
            end
            r_reg_prev <= 8'h00;
            g_reg_prev <= 8'h00;
            b_reg_prev <= 8'h00;
            frame_counter <= 8'h00;
        end else if (gx4000_mode) begin
            // Register writes
            if (cpu_wr) begin
                case (cpu_addr[7:0])
                    8'h80: screen_x <= cpu_data;
                    8'h81: screen_y <= cpu_data;
                    8'h82: video_mode <= cpu_data;
                    8'h83: collision_flags <= cpu_data;
                    
                    // Sprite transformation registers
                    8'h84: sprite_scale_x[cpu_addr[10:8]] <= cpu_data;
                    8'h85: sprite_scale_y[cpu_addr[10:8]] <= cpu_data;
                    8'h86: sprite_rotation[cpu_addr[10:8]] <= cpu_data;
                    8'h87: sprite_center_x[cpu_addr[10:8]] <= cpu_data;
                    8'h88: sprite_center_y[cpu_addr[10:8]] <= cpu_data;
                    8'h89: sprite_alpha[cpu_addr[10:8]] <= cpu_data;
                    8'h8A: sprite_flip_x[cpu_addr[10:8]] <= cpu_data;
                    8'h8B: sprite_flip_y[cpu_addr[10:8]] <= cpu_data;
                    8'h8C: sprite_priority[cpu_addr[10:8]] <= cpu_data;
                    8'h8D: sprite_effect[cpu_addr[10:8]] <= cpu_data;
                    
                    // Configuration registers
                    8'h90: config_mode <= cpu_data;
                    8'h91: config_palette <= cpu_data;
                    8'h92: config_sprite <= cpu_data;
                    8'h93: config_video <= cpu_data;
                    8'h94: config_audio <= cpu_data;
                    8'h95: config_io <= cpu_data;
                    
                    // Preset management
                    8'h96: config_preset <= cpu_data;
                    8'h97: config_save[cpu_addr[10:8]] <= cpu_data;
                    8'h98: config_load[cpu_addr[10:8]] <= cpu_data;
                endcase
                
                // Palette writes
                if (cpu_addr[15:8] == 8'h7F && cpu_addr[7:4] == 4'h6) begin
                    palette[cpu_addr[3:0]] <= {cpu_data, 16'h0000};
                end
            end
            
            // Video processing
            if (!hblank && !vblank) begin
                if (sprite_active) begin
                    // Get sprite transformation parameters
                    angle = sprite_rotation[active_sprite];
                    scale_x = sprite_scale_x[active_sprite];
                    scale_y = sprite_scale_y[active_sprite];
                    center_x = sprite_center_x[active_sprite];
                    center_y = sprite_center_y[active_sprite];
                    
                    // Apply scaling
                    rot_x = ((screen_x - center_x) * scale_x) >> 6;
                    rot_y = ((screen_y - center_y) * scale_y) >> 6;
                    
                    // Apply rotation
                    cos_angle = cos_table[angle];
                    sin_angle = sin_table[angle];
                    rot_x = (rot_x * cos_angle - rot_y * sin_angle) >> 8;
                    rot_y = (rot_x * sin_angle + rot_y * cos_angle) >> 8;
                    
                    // Apply flipping
                    if (sprite_flip_x[active_sprite]) begin
                        rot_x = -rot_x;
                    end
                    if (sprite_flip_y[active_sprite]) begin
                        rot_y = -rot_y;
                    end
                    
                    // Final position
                    final_x = center_x + rot_x[7:0];
                    final_y = center_y + rot_y[7:0];
                    
                    // Apply alpha blending
                    alpha = sprite_alpha[active_sprite];
                    r_reg <= (r_reg * alpha + r_reg_prev * (8'hFF - alpha)) >> 8;
                    g_reg <= (g_reg * alpha + g_reg_prev * (8'hFF - alpha)) >> 8;
                    b_reg <= (b_reg * alpha + b_reg_prev * (8'hFF - alpha)) >> 8;
                    
                    // Store previous values for effects
                    r_reg_prev <= r_reg;
                    g_reg_prev <= g_reg;
                    b_reg_prev <= b_reg;
                    
                    // Apply sprite effects
                    case (sprite_effect[active_sprite])
                        8'h00: begin // Normal
                            // No effect
                        end
                        8'h01: begin // Outline
                            if (sprite_pixel == 8'h00) begin
                                r_reg <= 8'hFF;
                                g_reg <= 8'hFF;
                                b_reg <= 8'hFF;
                            end
                        end
                        8'h02: begin // Shadow
                            r_reg <= r_reg >> 1;
                            g_reg <= g_reg >> 1;
                            b_reg <= b_reg >> 1;
                        end
                        8'h03: begin // Glow
                            r_reg <= (r_reg + 8'h80) >> 1;
                            g_reg <= (g_reg + 8'h80) >> 1;
                            b_reg <= (b_reg + 8'h80) >> 1;
                        end
                        8'h04: begin // Invert
                            r_reg <= ~r_reg;
                            g_reg <= ~g_reg;
                            b_reg <= ~b_reg;
                        end
                        8'h05: begin // Grayscale
                            gray = (r_reg + g_reg + b_reg) / 3;
                            r_reg <= gray;
                            g_reg <= gray;
                            b_reg <= gray;
                        end
                    endcase
                    
                    // Collision detection
                    if (collision_flags[sprite_id]) begin
                        collision_flags[sprite_id] <= 1'b0;
                    end
                end else begin
                    // Background color with video mode effects
                    case (video_mode)
                        8'h00: begin // Normal mode
                            r_reg <= palette[{r_in, 3'b000}][23:16];
                            g_reg <= palette[{g_in, 3'b000}][15:8];
                            b_reg <= palette[{b_in, 3'b000}][7:0];
                        end
                        8'h01: begin // Double width
                            r_reg <= palette[{r_in, 3'b000}][23:16];
                            g_reg <= palette[{g_in, 3'b000}][15:8];
                            b_reg <= palette[{b_in, 3'b000}][7:0];
                            if (screen_x[0]) begin
                                r_reg <= r_reg;
                                g_reg <= g_reg;
                                b_reg <= b_reg;
                            end
                        end
                        8'h02: begin // Double height
                            r_reg <= palette[{r_in, 3'b000}][23:16];
                            g_reg <= palette[{g_in, 3'b000}][15:8];
                            b_reg <= palette[{b_in, 3'b000}][7:0];
                            if (screen_y[0]) begin
                                r_reg <= r_reg;
                                g_reg <= g_reg;
                                b_reg <= b_reg;
                            end
                        end
                        8'h03: begin // Interlaced
                            r_reg <= palette[{r_in, 3'b000}][23:16];
                            g_reg <= palette[{g_in, 3'b000}][15:8];
                            b_reg <= palette[{b_in, 3'b000}][7:0];
                            if (screen_y[0]) begin
                                r_reg <= 8'h00;
                                g_reg <= 8'h00;
                                b_reg <= 8'h00;
                            end
                        end
                        8'h04: begin // Scanline
                            r_reg <= palette[{r_in, 3'b000}][23:16];
                            g_reg <= palette[{g_in, 3'b000}][15:8];
                            b_reg <= palette[{b_in, 3'b000}][7:0];
                            if (screen_y[0]) begin
                                r_reg <= r_reg >> 1;
                                g_reg <= g_reg >> 1;
                                b_reg <= b_reg >> 1;
                            end
                        end
                        8'h05: begin // Shadow
                            r_reg <= palette[{r_in, 3'b000}][23:16];
                            g_reg <= palette[{g_in, 3'b000}][15:8];
                            b_reg <= palette[{b_in, 3'b000}][7:0];
                            r_reg <= r_reg >> 1;
                            g_reg <= g_reg >> 1;
                            b_reg <= b_reg >> 1;
                        end
                        8'h06: begin // Ghost
                            r_reg <= palette[{r_in, 3'b000}][23:16];
                            g_reg <= palette[{g_in, 3'b000}][15:8];
                            b_reg <= palette[{b_in, 3'b000}][7:0];
                            r_reg <= (r_reg + 8'h80) >> 1;
                            g_reg <= (g_reg + 8'h80) >> 1;
                            b_reg <= (b_reg + 8'h80) >> 1;
                        end
                        8'h07: begin // Blur
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            r_reg <= (r_reg + r_reg_prev) >> 1;
                            g_reg <= (g_reg + g_reg_prev) >> 1;
                            b_reg <= (b_reg + b_reg_prev) >> 1;
                        end
                        8'h08: begin // Pixelate
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            if (screen_x[1:0] != 2'b00 || screen_y[1:0] != 2'b00) begin
                                r_reg <= r_reg_prev;
                                g_reg <= g_reg_prev;
                                b_reg <= b_reg_prev;
                            end
                        end
                        8'h09: begin // Wave
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            wave_offset = (screen_y * 8'h20) >> 8;
                            wave_x = screen_x + wave_offset;
                            if (wave_x[7:0] != screen_x[7:0]) begin
                                r_reg <= r_reg_prev;
                                g_reg <= g_reg_prev;
                                b_reg <= b_reg_prev;
                            end
                        end
                        8'h0A: begin // Zoom
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            zoom_x = (screen_x - 8'h40) * 8'h80 >> 7;
                            zoom_y = (screen_y - 8'h40) * 8'h80 >> 7;
                            if (zoom_x[7:0] != screen_x[7:0] || zoom_y[7:0] != screen_y[7:0]) begin
                                r_reg <= r_reg_prev;
                                g_reg <= g_reg_prev;
                                b_reg <= b_reg_prev;
                            end
                        end
                        8'h0B: begin // Color cycle
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            cycle_offset = (frame_counter * 8'h20) >> 8;
                            r_reg <= palette[(sprite_pixel[7:5] + cycle_offset) & 5'h1F][23:16];
                            g_reg <= palette[(sprite_pixel[4:2] + cycle_offset) & 5'h1F][15:8];
                            b_reg <= palette[(sprite_pixel[1:0] + cycle_offset) & 5'h1F][7:0];
                        end
                        8'h0C: begin // RGB shift
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            r_reg <= r_reg << 1;
                            g_reg <= g_reg >> 1;
                            b_reg <= b_reg << 1;
                        end
                        8'h0D: begin // CRT scanlines
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            if (screen_y[0]) begin
                                r_reg <= r_reg >> 2;
                                g_reg <= g_reg >> 2;
                                b_reg <= b_reg >> 2;
                            end
                        end
                        8'h0E: begin // CRT phosphor
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            r_reg <= (r_reg + (r_reg_prev >> 1)) >> 1;
                            g_reg <= (g_reg + (g_reg_prev >> 1)) >> 1;
                            b_reg <= (b_reg + (b_reg_prev >> 1)) >> 1;
                        end
                        8'h0F: begin // CRT bloom
                            r_reg <= palette[sprite_pixel[7:5]][23:16];
                            g_reg <= palette[sprite_pixel[4:2]][15:8];
                            b_reg <= palette[sprite_pixel[1:0]][7:0];
                            r_reg <= (r_reg + (r_reg_prev >> 2)) >> 1;
                            g_reg <= (g_reg + (g_reg_prev >> 2)) >> 1;
                            b_reg <= (b_reg + (b_reg_prev >> 2)) >> 1;
                        end
                    endcase
                end
            end
            
            // Apply configuration
            if (config_mode[0]) begin // Enable enhanced features
                // Apply palette configuration
                if (config_palette[0]) begin // Enable 32-color mode
                    // Use full 32-color palette
                end else begin
                    // Use 16-color mode
                    r_reg <= r_reg & 2'h3;
                    g_reg <= g_reg & 2'h3;
                    b_reg <= b_reg & 2'h3;
                end
                
                // Apply sprite configuration
                if (config_sprite[0]) begin // Enable sprite transformations
                    // Use transformed sprite coordinates
                end else begin
                    // Use original sprite coordinates
                end
                
                // Apply video configuration
                if (config_video[0]) begin // Enable video effects
                    // Use video mode effects
                end else begin
                    // Use normal video mode
                    video_mode <= 8'h00;
                end
                
                // Apply audio configuration
                if (config_audio[0]) begin // Enable enhanced audio
                    // Configure audio channels
                end
                
                // Apply I/O configuration
                if (config_io[0]) begin // Enable enhanced I/O
                    // Configure I/O ports
                end
                
                // Apply preset configuration
                if (config_preset[7]) begin // Load preset
                    case (config_preset[2:0])
                        3'h0: begin
                            config_mode <= config_load[0];
                            config_palette <= config_load[1];
                            config_sprite <= config_load[2];
                            config_video <= config_load[3];
                            config_audio <= config_load[4];
                            config_io <= config_load[5];
                        end
                        3'h1: begin
                            config_mode <= config_load[1];
                            config_palette <= config_load[2];
                            config_sprite <= config_load[3];
                            config_video <= config_load[4];
                            config_audio <= config_load[5];
                            config_io <= config_load[6];
                        end
                        // ... more preset cases ...
                    endcase
                end else if (config_preset[6]) begin // Save preset
                    case (config_preset[2:0])
                        3'h0: begin
                            config_save[0] <= config_mode;
                            config_save[1] <= config_palette;
                            config_save[2] <= config_sprite;
                            config_save[3] <= config_video;
                            config_save[4] <= config_audio;
                            config_save[5] <= config_io;
                        end
                        3'h1: begin
                            config_save[1] <= config_mode;
                            config_save[2] <= config_palette;
                            config_save[3] <= config_sprite;
                            config_save[4] <= config_video;
                            config_save[5] <= config_audio;
                            config_save[6] <= config_io;
                        end
                        // ... more preset cases ...
                    endcase
                end
            end else begin
                // Disable enhanced features
                video_mode <= 8'h00;
                r_reg <= 2'h0;
                g_reg <= 2'h0;
                b_reg <= 2'h0;
            end
            
            // Frame counter for effects
            if (vblank) begin
                frame_counter <= frame_counter + 1;
            end
        end
    end
    
    // Video output
    assign r_out = r_reg;
    assign g_out = g_reg;
    assign b_out = b_reg;
    
    // Collision register
    assign collision_reg = collision_flags;
    
    // Configuration register output
    assign config_reg = config_mode;

endmodule 